LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY dec3to8 IS
	PORT (w : IN STD_LOGIC_VECTOR(2 DOWNTO 0) ;
	y : OUT STD_LOGIC_VECTOR(0 TO 7) ) ;
END dec3to8 ;

ARCHITECTURE Behavior OF dec3to8 IS
BEGIN
	WITH w SELECT
		y <=  "10000000" WHEN "000",
				"01000000" WHEN "001",
				"00100000" WHEN "010",
				"00010000" WHEN "011",
				"00001000" WHEN "100",
				"00000100" WHEN "101",
				"00000010" WHEN "110",
				"00000001" WHEN "111",
				"00000000" WHEN OTHERS;
END Behavior ;